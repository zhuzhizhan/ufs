`timescale 1ns / 1ps
module Decode_8Bto10B(
	input	wire [9:0] data_in,
	input	wire       k_in,
	output	reg  [7:0] data_out
);
	        reg        rd_5bto6b;
	        reg  [4:0] lsb;
	        reg  [2:0] msb;
	        reg  [2:0] i;
                reg  [7:0] data_out;
			
    initial
		begin
			case(data_in[9:4])
				6'b100111:
					begin
						lsb=5'b00000;
						rd_5bto6b=1;
					end
				6'b011000:
					begin
						lsb=5'b00000;
						rd_5bto6b=0;
					end
				6'b011101:
					begin
						lsb=5'b00001;
						rd_5bto6b=1;
					end
				6'b100010:
					begin
						lsb=5'b00001;
						rd_5bto6b=0;
					end
				6'b101101:
					begin
						lsb=5'b00010;
						rd_5bto6b=1;
					end
				6'b010010:
					begin
						lsb=5'b00010;
						rd_5bto6b=0;
					end
				6'b110001:
					begin
						lsb=5'b00011;
						rd_5bto6b=0;
					end
				6'b110101:
					begin
						lsb=5'b00100;
						rd_5bto6b=1;
					end
				6'b001010:
					begin
						lsb=5'b00100;
						rd_5bto6b=0;
					end
				6'b101001:
					begin
						lsb=5'b00101;
						rd_5bto6b=0;
					end
				6'b011001:
					begin
						lsb=5'b00110;
						rd_5bto6b=0;
					end
				6'b111000:
					begin
						lsb=5'b00111;
						rd_5bto6b=1;
					end
				6'b000111:
					begin
						lsb=5'b00111;
						rd_5bto6b=1;
					end
				6'b111001:
					begin
						lsb=5'b01000;
						rd_5bto6b=1;
					end
				6'b000110:
					begin
						lsb=5'b01000;
						rd_5bto6b=0;
					end
				6'b100101:
					begin
						lsb=5'b01001;
						rd_5bto6b=0;
					end
				6'b010101:
					begin
						lsb=5'b01010;
						rd_5bto6b=0;
					end
				6'b110100:
					begin
						lsb=5'b01011;
						rd_5bto6b=1;
					end
				6'b001101:
					begin
						lsb=5'b01100;
						rd_5bto6b=0;
					end
				6'b101100:
					begin
						lsb=5'b01101;
						rd_5bto6b=1;
					end
				6'b011100:
					begin
						lsb=5'b01110;
						rd_5bto6b=1;
					end
				6'b010111:
					begin
						lsb=5'b01111;
						rd_5bto6b=1;
					end
				6'b101000:
					begin
						lsb=5'b01111;
						rd_5bto6b=0;
					end
				6'b011011:
					begin
						lsb=5'b10000;
						rd_5bto6b=1;
					end
				6'b100100:
					begin
						lsb=5'b10000;
						rd_5bto6b=0;
					end
				6'b100011:
					begin
						lsb=5'b10001;
						rd_5bto6b=0;
					end
				6'b010011:
					begin
						lsb=5'b10010;
						rd_5bto6b=0;
					end
				6'b110010:
					begin
						lsb=5'b10011;
						rd_5bto6b=1;
					end
				6'b001011:
					begin
						lsb=5'b10100;
						rd_5bto6b=0;
					end
				6'b101010:
					begin
						lsb=5'b10101;
						rd_5bto6b=1;
					end
				6'b011010:
					begin
						lsb=5'b10110;
						rd_5bto6b=1;
					end
				6'b111010:
					begin
						lsb=5'b10111;
						rd_5bto6b=1;
					end
				6'b000101:
					begin
						lsb=5'b10111;
						rd_5bto6b=0;
					end
				6'b110011:
					begin
						lsb=5'b11000;
						rd_5bto6b=1;
					end
				6'b001100:
					begin
						lsb=5'b11000;
						rd_5bto6b=0;
					end
				6'b100110:
					begin
						lsb=5'b11001;
					   rd_5bto6b=1;
					end
				6'b010110:
					begin
						lsb=5'b11010;
						rd_5bto6b=1;
					end
				6'b110110:
					begin
						lsb=5'b11011;
						rd_5bto6b=1;
					end
				6'b001001:
					begin
						lsb=5'b11011;
						rd_5bto6b=0;
					end
				6'b001110:
					begin
						lsb=5'b11100;
						rd_5bto6b=1;
					end
				6'b101110:
					begin
						lsb=5'b11101;
						rd_5bto6b=1;
					end
				6'b010001:
					begin
						lsb=5'b11101;
						rd_5bto6b=0;
					end
				6'b011110:
					begin
						lsb=5'b11110;
						rd_5bto6b=1;
					end
				6'b100001:
					begin
						lsb=5'b11110;
						rd_5bto6b=0;
					end
				6'b101011:
					begin
						lsb=5'b11111;
						rd_5bto6b=1;
					end
				6'b010100:
					begin
						lsb=5'b11111;
						rd_5bto6b=0;
					end
				6'b001111:
					begin
						lsb=5'b11100;
						rd_5bto6b=1;
					end
				6'b110000:
					begin
						lsb=5'b11100;
						rd_5bto6b=0;
					end
				default:
					begin
						lsb=5'bXXXXX;
						rd_5bto6b=1'bX;
					end
		 endcase
		 
		for(i=0;i<5;i=i+1)
			data_out[i]=lsb[i];
			
	    if(k_in)
			begin
				if(rd_5bto6b)
					case(data_in[3:0])
						4'b0100:
							msb=3'b000;
						4'b1001:
							msb=3'b001;
						4'b0101:
							msb=3'b010;
						4'b0011:
							msb=3'b011;
						4'b0010:
							msb=3'b100;
						4'b1010:
							msb=3'b101;
						4'b0110:
							msb=3'b110;
						4'b1000:
							msb=3'b111;
						default:
							msb=3'bXXX;
					endcase
				else
					case(data_in[3:0])
						4'b1011:
							msb=3'b000;
						4'b0110:
							msb=3'b001;
						4'b1010:
							msb=3'b010;
						4'b1100:
							msb=3'b011;
						4'b1101:
							msb=3'b100;
						4'b0101:
							msb=3'b101;
						4'b1001:
							msb=3'b110;
						4'b0111:
							msb=3'b111;
						default:
							msb=3'bXXX;
					endcase
			end
		else
			begin
				if(rd_5bto6b)
					case(data_in[3:0])
						4'b0100:
							msb=3'b000;
						4'b1001:
							msb=3'b001;
						4'b0101:
							msb=3'b010;
						4'b0011:
							msb=3'b011;
						4'b0010:
							msb=3'b100;
						4'b1010:
							msb=3'b101;
						4'b0110:
							msb=3'b110;
						4'b0001:
							msb=3'b111;
						4'b1000:
							msb=3'b111;
						default:
							msb=3'bXXX;
					endcase
				else
					case(data_in[3:0])
						4'b1011:
							msb=3'b000;
						4'b1001:
							msb=3'b001;
						4'b0101:
							msb=3'b010;
						4'b1100:
							msb=3'b011;
						4'b1101:
							msb=3'b100;
						4'b1010:
							msb=3'b101;
						4'b0110:
							msb=3'b110;
						4'b1110:
							msb=3'b111;
						4'b0111:
							msb=3'b111;
						default:
							msb=3'bXXX;
					endcase
			end
				
		   
			for(i=0;i<3;i=i+1)
				data_out[i+5]=msb[i];
				
		end
		
endmodule



module testbench;

	reg  [9:0] data_in;
	reg        k_in;
	wire [7:0] data_out;
	
	Decode_8Bto10B  testbench(.data_in(),.k_in(k_in),.data_out(data_out));
	
	initial 
		begin
			data_in=10'b1100001001;
			k_in=0;
		end
	
endmodule
